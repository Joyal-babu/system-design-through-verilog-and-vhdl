library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity fa is
    Port (
           A    : in  STD_LOGIC;
           B    : in  STD_LOGIC;
           Cin  : in  STD_LOGIC;
           Sum  : out STD_LOGIC;
           Cout : out STD_LOGIC );
end fa;

architecture Behavioral of fa is

begin
    Sum  <= (A xor B xor Cin);
    Cout <= (A and B) or (B and Cin) or (A and Cin);

end Behavioral;
